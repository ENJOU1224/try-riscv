/* 
    -- ============================================================================
    -- FILE NAME	: decode.v
    -- DESCRIPTION : 指令集架构
    -- ----------------------------------------------------------------------------
    -- Revision  Date		  Coding_by	 Comment
    -- 1.0.0	  2021/09/28  enjou		 初版
    -- ============================================================================
*/

module decode (
    input   [63:0]  i_PC_64,
    input   [31:0]  i_Inst_32,
    input   [63:0]  i_GRFData1_64,
    input   [63:0]  i_GRFData2_64,
    input   [63:0]  i_CSRData_64,
);
endmodule